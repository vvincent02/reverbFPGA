// reverbFPGA_Qsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module reverbFPGA_Qsys (
		input  wire  clk_clk  // clk.clk
	);

	wire    hps_0_h2f_reset_reset;          // hps_0:h2f_rst_n -> rst_controller:reset_in0
	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> pio_0:reset_n

	reverbFPGA_Qsys_hps_0 #(
		.F2S_Width (1),
		.S2F_Width (1)
	) hps_0 (
		.h2f_mpu_eventi     (),                      //    h2f_mpu_events.eventi
		.h2f_mpu_evento     (),                      //                  .evento
		.h2f_mpu_standbywfe (),                      //                  .standbywfe
		.h2f_mpu_standbywfi (),                      //                  .standbywfi
		.mem_a              (),                      //            memory.mem_a
		.mem_ba             (),                      //                  .mem_ba
		.mem_ck             (),                      //                  .mem_ck
		.mem_ck_n           (),                      //                  .mem_ck_n
		.mem_cke            (),                      //                  .mem_cke
		.mem_cs_n           (),                      //                  .mem_cs_n
		.mem_ras_n          (),                      //                  .mem_ras_n
		.mem_cas_n          (),                      //                  .mem_cas_n
		.mem_we_n           (),                      //                  .mem_we_n
		.mem_reset_n        (),                      //                  .mem_reset_n
		.mem_dq             (),                      //                  .mem_dq
		.mem_dqs            (),                      //                  .mem_dqs
		.mem_dqs_n          (),                      //                  .mem_dqs_n
		.mem_odt            (),                      //                  .mem_odt
		.mem_dm             (),                      //                  .mem_dm
		.oct_rzqin          (),                      //                  .oct_rzqin
		.h2f_rst_n          (hps_0_h2f_reset_reset), //         h2f_reset.reset_n
		.f2h_sdram0_clk     (clk_clk),               //  f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR  (),                      //   f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN   (),                      //                  .arlen
		.f2h_sdram0_ARID    (),                      //                  .arid
		.f2h_sdram0_ARSIZE  (),                      //                  .arsize
		.f2h_sdram0_ARBURST (),                      //                  .arburst
		.f2h_sdram0_ARLOCK  (),                      //                  .arlock
		.f2h_sdram0_ARPROT  (),                      //                  .arprot
		.f2h_sdram0_ARVALID (),                      //                  .arvalid
		.f2h_sdram0_ARCACHE (),                      //                  .arcache
		.f2h_sdram0_AWADDR  (),                      //                  .awaddr
		.f2h_sdram0_AWLEN   (),                      //                  .awlen
		.f2h_sdram0_AWID    (),                      //                  .awid
		.f2h_sdram0_AWSIZE  (),                      //                  .awsize
		.f2h_sdram0_AWBURST (),                      //                  .awburst
		.f2h_sdram0_AWLOCK  (),                      //                  .awlock
		.f2h_sdram0_AWPROT  (),                      //                  .awprot
		.f2h_sdram0_AWVALID (),                      //                  .awvalid
		.f2h_sdram0_AWCACHE (),                      //                  .awcache
		.f2h_sdram0_BRESP   (),                      //                  .bresp
		.f2h_sdram0_BID     (),                      //                  .bid
		.f2h_sdram0_BVALID  (),                      //                  .bvalid
		.f2h_sdram0_BREADY  (),                      //                  .bready
		.f2h_sdram0_ARREADY (),                      //                  .arready
		.f2h_sdram0_AWREADY (),                      //                  .awready
		.f2h_sdram0_RREADY  (),                      //                  .rready
		.f2h_sdram0_RDATA   (),                      //                  .rdata
		.f2h_sdram0_RRESP   (),                      //                  .rresp
		.f2h_sdram0_RLAST   (),                      //                  .rlast
		.f2h_sdram0_RID     (),                      //                  .rid
		.f2h_sdram0_RVALID  (),                      //                  .rvalid
		.f2h_sdram0_WLAST   (),                      //                  .wlast
		.f2h_sdram0_WVALID  (),                      //                  .wvalid
		.f2h_sdram0_WDATA   (),                      //                  .wdata
		.f2h_sdram0_WSTRB   (),                      //                  .wstrb
		.f2h_sdram0_WREADY  (),                      //                  .wready
		.f2h_sdram0_WID     (),                      //                  .wid
		.h2f_axi_clk        (clk_clk),               //     h2f_axi_clock.clk
		.h2f_AWID           (),                      //    h2f_axi_master.awid
		.h2f_AWADDR         (),                      //                  .awaddr
		.h2f_AWLEN          (),                      //                  .awlen
		.h2f_AWSIZE         (),                      //                  .awsize
		.h2f_AWBURST        (),                      //                  .awburst
		.h2f_AWLOCK         (),                      //                  .awlock
		.h2f_AWCACHE        (),                      //                  .awcache
		.h2f_AWPROT         (),                      //                  .awprot
		.h2f_AWVALID        (),                      //                  .awvalid
		.h2f_AWREADY        (),                      //                  .awready
		.h2f_WID            (),                      //                  .wid
		.h2f_WDATA          (),                      //                  .wdata
		.h2f_WSTRB          (),                      //                  .wstrb
		.h2f_WLAST          (),                      //                  .wlast
		.h2f_WVALID         (),                      //                  .wvalid
		.h2f_WREADY         (),                      //                  .wready
		.h2f_BID            (),                      //                  .bid
		.h2f_BRESP          (),                      //                  .bresp
		.h2f_BVALID         (),                      //                  .bvalid
		.h2f_BREADY         (),                      //                  .bready
		.h2f_ARID           (),                      //                  .arid
		.h2f_ARADDR         (),                      //                  .araddr
		.h2f_ARLEN          (),                      //                  .arlen
		.h2f_ARSIZE         (),                      //                  .arsize
		.h2f_ARBURST        (),                      //                  .arburst
		.h2f_ARLOCK         (),                      //                  .arlock
		.h2f_ARCACHE        (),                      //                  .arcache
		.h2f_ARPROT         (),                      //                  .arprot
		.h2f_ARVALID        (),                      //                  .arvalid
		.h2f_ARREADY        (),                      //                  .arready
		.h2f_RID            (),                      //                  .rid
		.h2f_RDATA          (),                      //                  .rdata
		.h2f_RRESP          (),                      //                  .rresp
		.h2f_RLAST          (),                      //                  .rlast
		.h2f_RVALID         (),                      //                  .rvalid
		.h2f_RREADY         (),                      //                  .rready
		.f2h_axi_clk        (clk_clk),               //     f2h_axi_clock.clk
		.f2h_AWID           (),                      //     f2h_axi_slave.awid
		.f2h_AWADDR         (),                      //                  .awaddr
		.f2h_AWLEN          (),                      //                  .awlen
		.f2h_AWSIZE         (),                      //                  .awsize
		.f2h_AWBURST        (),                      //                  .awburst
		.f2h_AWLOCK         (),                      //                  .awlock
		.f2h_AWCACHE        (),                      //                  .awcache
		.f2h_AWPROT         (),                      //                  .awprot
		.f2h_AWVALID        (),                      //                  .awvalid
		.f2h_AWREADY        (),                      //                  .awready
		.f2h_AWUSER         (),                      //                  .awuser
		.f2h_WID            (),                      //                  .wid
		.f2h_WDATA          (),                      //                  .wdata
		.f2h_WSTRB          (),                      //                  .wstrb
		.f2h_WLAST          (),                      //                  .wlast
		.f2h_WVALID         (),                      //                  .wvalid
		.f2h_WREADY         (),                      //                  .wready
		.f2h_BID            (),                      //                  .bid
		.f2h_BRESP          (),                      //                  .bresp
		.f2h_BVALID         (),                      //                  .bvalid
		.f2h_BREADY         (),                      //                  .bready
		.f2h_ARID           (),                      //                  .arid
		.f2h_ARADDR         (),                      //                  .araddr
		.f2h_ARLEN          (),                      //                  .arlen
		.f2h_ARSIZE         (),                      //                  .arsize
		.f2h_ARBURST        (),                      //                  .arburst
		.f2h_ARLOCK         (),                      //                  .arlock
		.f2h_ARCACHE        (),                      //                  .arcache
		.f2h_ARPROT         (),                      //                  .arprot
		.f2h_ARVALID        (),                      //                  .arvalid
		.f2h_ARREADY        (),                      //                  .arready
		.f2h_ARUSER         (),                      //                  .aruser
		.f2h_RID            (),                      //                  .rid
		.f2h_RDATA          (),                      //                  .rdata
		.f2h_RRESP          (),                      //                  .rresp
		.f2h_RLAST          (),                      //                  .rlast
		.f2h_RVALID         (),                      //                  .rvalid
		.f2h_RREADY         (),                      //                  .rready
		.h2f_lw_axi_clk     (clk_clk),               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID        (),                      // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR      (),                      //                  .awaddr
		.h2f_lw_AWLEN       (),                      //                  .awlen
		.h2f_lw_AWSIZE      (),                      //                  .awsize
		.h2f_lw_AWBURST     (),                      //                  .awburst
		.h2f_lw_AWLOCK      (),                      //                  .awlock
		.h2f_lw_AWCACHE     (),                      //                  .awcache
		.h2f_lw_AWPROT      (),                      //                  .awprot
		.h2f_lw_AWVALID     (),                      //                  .awvalid
		.h2f_lw_AWREADY     (),                      //                  .awready
		.h2f_lw_WID         (),                      //                  .wid
		.h2f_lw_WDATA       (),                      //                  .wdata
		.h2f_lw_WSTRB       (),                      //                  .wstrb
		.h2f_lw_WLAST       (),                      //                  .wlast
		.h2f_lw_WVALID      (),                      //                  .wvalid
		.h2f_lw_WREADY      (),                      //                  .wready
		.h2f_lw_BID         (),                      //                  .bid
		.h2f_lw_BRESP       (),                      //                  .bresp
		.h2f_lw_BVALID      (),                      //                  .bvalid
		.h2f_lw_BREADY      (),                      //                  .bready
		.h2f_lw_ARID        (),                      //                  .arid
		.h2f_lw_ARADDR      (),                      //                  .araddr
		.h2f_lw_ARLEN       (),                      //                  .arlen
		.h2f_lw_ARSIZE      (),                      //                  .arsize
		.h2f_lw_ARBURST     (),                      //                  .arburst
		.h2f_lw_ARLOCK      (),                      //                  .arlock
		.h2f_lw_ARCACHE     (),                      //                  .arcache
		.h2f_lw_ARPROT      (),                      //                  .arprot
		.h2f_lw_ARVALID     (),                      //                  .arvalid
		.h2f_lw_ARREADY     (),                      //                  .arready
		.h2f_lw_RID         (),                      //                  .rid
		.h2f_lw_RDATA       (),                      //                  .rdata
		.h2f_lw_RRESP       (),                      //                  .rresp
		.h2f_lw_RLAST       (),                      //                  .rlast
		.h2f_lw_RVALID      (),                      //                  .rvalid
		.h2f_lw_RREADY      ()                       //                  .rready
	);

	reverbFPGA_Qsys_pio_0 pio_0 (
		.clk        (clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset), //               reset.reset_n
		.address    (),                                //                  s1.address
		.write_n    (),                                //                    .write_n
		.writedata  (),                                //                    .writedata
		.chipselect (),                                //                    .chipselect
		.readdata   (),                                //                    .readdata
		.bidir_port ()                                 // external_connection.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
