-- altclkctrl_inst.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity altclkctrl_inst is
	port (
		inclk  : in  std_logic := '0'; --  altclkctrl_input.inclk
		ena    : in  std_logic := '0'; --                  .ena
		outclk : out std_logic         -- altclkctrl_output.outclk
	);
end entity altclkctrl_inst;

architecture rtl of altclkctrl_inst is
	component reverbFPGA_Qsys_serial_flash_loader_altclkctrl_inst_altclkctrl_inst is
		port (
			inclk  : in  std_logic := 'X'; -- inclk
			ena    : in  std_logic := 'X'; -- ena
			outclk : out std_logic         -- outclk
		);
	end component reverbFPGA_Qsys_serial_flash_loader_altclkctrl_inst_altclkctrl_inst;

begin

	altclkctrl_inst : component reverbFPGA_Qsys_serial_flash_loader_altclkctrl_inst_altclkctrl_inst
		port map (
			inclk  => inclk,  --  altclkctrl_input.inclk
			ena    => ena,    --                  .ena
			outclk => outclk  -- altclkctrl_output.outclk
		);

end architecture rtl; -- of altclkctrl_inst
