-- reverbFPGA_Qsys.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity reverbFPGA_Qsys is
	port (
		audio_controller_avalon_left_channel_sink_data     : in    std_logic_vector(23 downto 0) := (others => '0'); --    audio_controller_avalon_left_channel_sink.data
		audio_controller_avalon_left_channel_sink_valid    : in    std_logic                     := '0';             --                                             .valid
		audio_controller_avalon_left_channel_sink_ready    : out   std_logic;                                        --                                             .ready
		audio_controller_avalon_left_channel_source_ready  : in    std_logic                     := '0';             --  audio_controller_avalon_left_channel_source.ready
		audio_controller_avalon_left_channel_source_data   : out   std_logic_vector(23 downto 0);                    --                                             .data
		audio_controller_avalon_left_channel_source_valid  : out   std_logic;                                        --                                             .valid
		audio_controller_avalon_right_channel_sink_data    : in    std_logic_vector(23 downto 0) := (others => '0'); --   audio_controller_avalon_right_channel_sink.data
		audio_controller_avalon_right_channel_sink_valid   : in    std_logic                     := '0';             --                                             .valid
		audio_controller_avalon_right_channel_sink_ready   : out   std_logic;                                        --                                             .ready
		audio_controller_avalon_right_channel_source_ready : in    std_logic                     := '0';             -- audio_controller_avalon_right_channel_source.ready
		audio_controller_avalon_right_channel_source_data  : out   std_logic_vector(23 downto 0);                    --                                             .data
		audio_controller_avalon_right_channel_source_valid : out   std_logic;                                        --                                             .valid
		audio_controller_external_interface_ADCDAT         : in    std_logic                     := '0';             --          audio_controller_external_interface.ADCDAT
		audio_controller_external_interface_ADCLRCK        : in    std_logic                     := '0';             --                                             .ADCLRCK
		audio_controller_external_interface_BCLK           : in    std_logic                     := '0';             --                                             .BCLK
		audio_controller_external_interface_DACDAT         : out   std_logic;                                        --                                             .DACDAT
		audio_controller_external_interface_DACLRCK        : in    std_logic                     := '0';             --                                             .DACLRCK
		audio_pll_0_audio_clk_clk                          : out   std_logic;                                        --                        audio_pll_0_audio_clk.clk
		clk_clk                                            : in    std_logic                     := '0';             --                                          clk.clk
		clksampling_clk                                    : out   std_logic;                                        --                                  clksampling.clk
		hps_0_h2f_mpu_events_eventi                        : in    std_logic                     := '0';             --                         hps_0_h2f_mpu_events.eventi
		hps_0_h2f_mpu_events_evento                        : out   std_logic;                                        --                                             .evento
		hps_0_h2f_mpu_events_standbywfe                    : out   std_logic_vector(1 downto 0);                     --                                             .standbywfe
		hps_0_h2f_mpu_events_standbywfi                    : out   std_logic_vector(1 downto 0);                     --                                             .standbywfi
		hps_io_hps_io_uart0_inst_RX                        : in    std_logic                     := '0';             --                                       hps_io.hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX                        : out   std_logic;                                        --                                             .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c1_inst_SDA                        : inout std_logic                     := '0';             --                                             .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL                        : inout std_logic                     := '0';             --                                             .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO48                     : inout std_logic                     := '0';             --                                             .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO53                     : inout std_logic                     := '0';             --                                             .hps_io_gpio_inst_GPIO53
		memory_mem_a                                       : out   std_logic_vector(14 downto 0);                    --                                       memory.mem_a
		memory_mem_ba                                      : out   std_logic_vector(2 downto 0);                     --                                             .mem_ba
		memory_mem_ck                                      : out   std_logic;                                        --                                             .mem_ck
		memory_mem_ck_n                                    : out   std_logic;                                        --                                             .mem_ck_n
		memory_mem_cke                                     : out   std_logic;                                        --                                             .mem_cke
		memory_mem_cs_n                                    : out   std_logic;                                        --                                             .mem_cs_n
		memory_mem_ras_n                                   : out   std_logic;                                        --                                             .mem_ras_n
		memory_mem_cas_n                                   : out   std_logic;                                        --                                             .mem_cas_n
		memory_mem_we_n                                    : out   std_logic;                                        --                                             .mem_we_n
		memory_mem_reset_n                                 : out   std_logic;                                        --                                             .mem_reset_n
		memory_mem_dq                                      : inout std_logic_vector(31 downto 0) := (others => '0'); --                                             .mem_dq
		memory_mem_dqs                                     : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                             .mem_dqs
		memory_mem_dqs_n                                   : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                             .mem_dqs_n
		memory_mem_odt                                     : out   std_logic;                                        --                                             .mem_odt
		memory_mem_dm                                      : out   std_logic_vector(3 downto 0);                     --                                             .mem_dm
		memory_oct_rzqin                                   : in    std_logic                     := '0';             --                                             .oct_rzqin
		reset_reset_n                                      : in    std_logic                     := '0';             --                                        reset.reset_n
		serial_flash_loader_0_noe_in_noe                   : in    std_logic                     := '0'              --                 serial_flash_loader_0_noe_in.noe
	);
end entity reverbFPGA_Qsys;

architecture rtl of reverbFPGA_Qsys is
	component reverbFPGA_Qsys_audio_controller is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset                        : in  std_logic                     := 'X';             -- reset
			from_adc_left_channel_ready  : in  std_logic                     := 'X';             -- ready
			from_adc_left_channel_data   : out std_logic_vector(23 downto 0);                    -- data
			from_adc_left_channel_valid  : out std_logic;                                        -- valid
			from_adc_right_channel_ready : in  std_logic                     := 'X';             -- ready
			from_adc_right_channel_data  : out std_logic_vector(23 downto 0);                    -- data
			from_adc_right_channel_valid : out std_logic;                                        -- valid
			to_dac_left_channel_data     : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_left_channel_valid    : in  std_logic                     := 'X';             -- valid
			to_dac_left_channel_ready    : out std_logic;                                        -- ready
			to_dac_right_channel_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_right_channel_valid   : in  std_logic                     := 'X';             -- valid
			to_dac_right_channel_ready   : out std_logic;                                        -- ready
			AUD_ADCDAT                   : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK                  : in  std_logic                     := 'X';             -- export
			AUD_BCLK                     : in  std_logic                     := 'X';             -- export
			AUD_DACDAT                   : out std_logic;                                        -- export
			AUD_DACLRCK                  : in  std_logic                     := 'X'              -- export
		);
	end component reverbFPGA_Qsys_audio_controller;

	component reverbFPGA_Qsys_audio_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component reverbFPGA_Qsys_audio_pll_0;

	component reverbFPGA_Qsys_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_mpu_eventi          : in    std_logic                     := 'X';             -- eventi
			h2f_mpu_evento          : out   std_logic;                                        -- evento
			h2f_mpu_standbywfe      : out   std_logic_vector(1 downto 0);                     -- standbywfe
			h2f_mpu_standbywfi      : out   std_logic_vector(1 downto 0);                     -- standbywfi
			mem_a                   : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                  : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                  : out   std_logic;                                        -- mem_ck
			mem_ck_n                : out   std_logic;                                        -- mem_ck_n
			mem_cke                 : out   std_logic;                                        -- mem_cke
			mem_cs_n                : out   std_logic;                                        -- mem_cs_n
			mem_ras_n               : out   std_logic;                                        -- mem_ras_n
			mem_cas_n               : out   std_logic;                                        -- mem_cas_n
			mem_we_n                : out   std_logic;                                        -- mem_we_n
			mem_reset_n             : out   std_logic;                                        -- mem_reset_n
			mem_dq                  : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                 : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n               : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                 : out   std_logic;                                        -- mem_odt
			mem_dm                  : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin               : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_uart0_inst_RX    : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX    : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c1_inst_SDA    : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL    : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO48 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			h2f_rst_n               : out   std_logic;                                        -- reset_n
			h2f_axi_clk             : in    std_logic                     := 'X';             -- clk
			h2f_AWID                : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR              : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN               : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE              : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST             : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK              : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE             : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT              : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID             : out   std_logic;                                        -- awvalid
			h2f_AWREADY             : in    std_logic                     := 'X';             -- awready
			h2f_WID                 : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA               : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_WSTRB               : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_WLAST               : out   std_logic;                                        -- wlast
			h2f_WVALID              : out   std_logic;                                        -- wvalid
			h2f_WREADY              : in    std_logic                     := 'X';             -- wready
			h2f_BID                 : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID              : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY              : out   std_logic;                                        -- bready
			h2f_ARID                : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR              : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN               : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE              : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST             : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK              : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE             : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT              : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID             : out   std_logic;                                        -- arvalid
			h2f_ARREADY             : in    std_logic                     := 'X';             -- arready
			h2f_RID                 : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST               : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID              : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY              : out   std_logic;                                        -- rready
			f2h_axi_clk             : in    std_logic                     := 'X';             -- clk
			f2h_AWID                : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- awid
			f2h_AWADDR              : in    std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			f2h_AWLEN               : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			f2h_AWSIZE              : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			f2h_AWBURST             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			f2h_AWLOCK              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			f2h_AWCACHE             : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			f2h_AWPROT              : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			f2h_AWVALID             : in    std_logic                     := 'X';             -- awvalid
			f2h_AWREADY             : out   std_logic;                                        -- awready
			f2h_AWUSER              : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- awuser
			f2h_WID                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wid
			f2h_WDATA               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB               : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST               : in    std_logic                     := 'X';             -- wlast
			f2h_WVALID              : in    std_logic                     := 'X';             -- wvalid
			f2h_WREADY              : out   std_logic;                                        -- wready
			f2h_BID                 : out   std_logic_vector(7 downto 0);                     -- bid
			f2h_BRESP               : out   std_logic_vector(1 downto 0);                     -- bresp
			f2h_BVALID              : out   std_logic;                                        -- bvalid
			f2h_BREADY              : in    std_logic                     := 'X';             -- bready
			f2h_ARID                : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- arid
			f2h_ARADDR              : in    std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			f2h_ARLEN               : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			f2h_ARSIZE              : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			f2h_ARBURST             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			f2h_ARLOCK              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			f2h_ARCACHE             : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			f2h_ARPROT              : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			f2h_ARVALID             : in    std_logic                     := 'X';             -- arvalid
			f2h_ARREADY             : out   std_logic;                                        -- arready
			f2h_ARUSER              : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- aruser
			f2h_RID                 : out   std_logic_vector(7 downto 0);                     -- rid
			f2h_RDATA               : out   std_logic_vector(31 downto 0);                    -- rdata
			f2h_RRESP               : out   std_logic_vector(1 downto 0);                     -- rresp
			f2h_RLAST               : out   std_logic;                                        -- rlast
			f2h_RVALID              : out   std_logic;                                        -- rvalid
			f2h_RREADY              : in    std_logic                     := 'X';             -- rready
			h2f_lw_axi_clk          : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID             : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR           : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN            : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE           : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST          : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK           : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE          : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT           : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID          : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY          : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID              : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA            : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB            : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST            : out   std_logic;                                        -- wlast
			h2f_lw_WVALID           : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY           : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID              : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP            : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID           : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY           : out   std_logic;                                        -- bready
			h2f_lw_ARID             : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR           : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN            : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE           : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST          : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK           : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE          : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT           : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID          : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY          : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID              : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA            : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP            : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST            : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID           : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY           : out   std_logic                                         -- rready
		);
	end component reverbFPGA_Qsys_hps_0;

	component altera_serial_flash_loader is
		generic (
			INTENDED_DEVICE_FAMILY  : string  := "";
			ENHANCED_MODE           : boolean := true;
			ENABLE_SHARED_ACCESS    : string  := "OFF";
			ENABLE_QUAD_SPI_SUPPORT : boolean := false;
			NCSO_WIDTH              : integer := 1
		);
		port (
			noe_in : in std_logic := 'X'  -- noe
		);
	end component altera_serial_flash_loader;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal rst_controller_reset_out_reset : std_logic; -- rst_controller:reset_out -> audio_controller:reset
	signal reset_reset_n_ports_inv        : std_logic; -- reset_reset_n:inv -> [audio_pll_0:ref_reset_reset, rst_controller:reset_in0]

begin

	audio_controller : component reverbFPGA_Qsys_audio_controller
		port map (
			clk                          => clk_clk,                                            --                         clk.clk
			reset                        => rst_controller_reset_out_reset,                     --                       reset.reset
			from_adc_left_channel_ready  => audio_controller_avalon_left_channel_source_ready,  --  avalon_left_channel_source.ready
			from_adc_left_channel_data   => audio_controller_avalon_left_channel_source_data,   --                            .data
			from_adc_left_channel_valid  => audio_controller_avalon_left_channel_source_valid,  --                            .valid
			from_adc_right_channel_ready => audio_controller_avalon_right_channel_source_ready, -- avalon_right_channel_source.ready
			from_adc_right_channel_data  => audio_controller_avalon_right_channel_source_data,  --                            .data
			from_adc_right_channel_valid => audio_controller_avalon_right_channel_source_valid, --                            .valid
			to_dac_left_channel_data     => audio_controller_avalon_left_channel_sink_data,     --    avalon_left_channel_sink.data
			to_dac_left_channel_valid    => audio_controller_avalon_left_channel_sink_valid,    --                            .valid
			to_dac_left_channel_ready    => audio_controller_avalon_left_channel_sink_ready,    --                            .ready
			to_dac_right_channel_data    => audio_controller_avalon_right_channel_sink_data,    --   avalon_right_channel_sink.data
			to_dac_right_channel_valid   => audio_controller_avalon_right_channel_sink_valid,   --                            .valid
			to_dac_right_channel_ready   => audio_controller_avalon_right_channel_sink_ready,   --                            .ready
			AUD_ADCDAT                   => audio_controller_external_interface_ADCDAT,         --          external_interface.export
			AUD_ADCLRCK                  => audio_controller_external_interface_ADCLRCK,        --                            .export
			AUD_BCLK                     => audio_controller_external_interface_BCLK,           --                            .export
			AUD_DACDAT                   => audio_controller_external_interface_DACDAT,         --                            .export
			AUD_DACLRCK                  => audio_controller_external_interface_DACLRCK         --                            .export
		);

	audio_pll_0 : component reverbFPGA_Qsys_audio_pll_0
		port map (
			ref_clk_clk        => clk_clk,                   --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,   --    ref_reset.reset
			audio_clk_clk      => audio_pll_0_audio_clk_clk, --    audio_clk.clk
			reset_source_reset => open                       -- reset_source.reset
		);

	hps_0 : component reverbFPGA_Qsys_hps_0
		generic map (
			F2S_Width => 1,
			S2F_Width => 1
		)
		port map (
			h2f_mpu_eventi          => hps_0_h2f_mpu_events_eventi,     --    h2f_mpu_events.eventi
			h2f_mpu_evento          => hps_0_h2f_mpu_events_evento,     --                  .evento
			h2f_mpu_standbywfe      => hps_0_h2f_mpu_events_standbywfe, --                  .standbywfe
			h2f_mpu_standbywfi      => hps_0_h2f_mpu_events_standbywfi, --                  .standbywfi
			mem_a                   => memory_mem_a,                    --            memory.mem_a
			mem_ba                  => memory_mem_ba,                   --                  .mem_ba
			mem_ck                  => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n                => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                 => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n                => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n               => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n               => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n             => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq                  => memory_mem_dq,                   --                  .mem_dq
			mem_dqs                 => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n               => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                 => memory_mem_odt,                  --                  .mem_odt
			mem_dm                  => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin               => memory_oct_rzqin,                --                  .oct_rzqin
			hps_io_uart0_inst_RX    => hps_io_hps_io_uart0_inst_RX,     --            hps_io.hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX    => hps_io_hps_io_uart0_inst_TX,     --                  .hps_io_uart0_inst_TX
			hps_io_i2c1_inst_SDA    => hps_io_hps_io_i2c1_inst_SDA,     --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL    => hps_io_hps_io_i2c1_inst_SCL,     --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO48 => hps_io_hps_io_gpio_inst_GPIO48,  --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53 => hps_io_hps_io_gpio_inst_GPIO53,  --                  .hps_io_gpio_inst_GPIO53
			h2f_rst_n               => open,                            --         h2f_reset.reset_n
			h2f_axi_clk             => clk_clk,                         --     h2f_axi_clock.clk
			h2f_AWID                => open,                            --    h2f_axi_master.awid
			h2f_AWADDR              => open,                            --                  .awaddr
			h2f_AWLEN               => open,                            --                  .awlen
			h2f_AWSIZE              => open,                            --                  .awsize
			h2f_AWBURST             => open,                            --                  .awburst
			h2f_AWLOCK              => open,                            --                  .awlock
			h2f_AWCACHE             => open,                            --                  .awcache
			h2f_AWPROT              => open,                            --                  .awprot
			h2f_AWVALID             => open,                            --                  .awvalid
			h2f_AWREADY             => open,                            --                  .awready
			h2f_WID                 => open,                            --                  .wid
			h2f_WDATA               => open,                            --                  .wdata
			h2f_WSTRB               => open,                            --                  .wstrb
			h2f_WLAST               => open,                            --                  .wlast
			h2f_WVALID              => open,                            --                  .wvalid
			h2f_WREADY              => open,                            --                  .wready
			h2f_BID                 => open,                            --                  .bid
			h2f_BRESP               => open,                            --                  .bresp
			h2f_BVALID              => open,                            --                  .bvalid
			h2f_BREADY              => open,                            --                  .bready
			h2f_ARID                => open,                            --                  .arid
			h2f_ARADDR              => open,                            --                  .araddr
			h2f_ARLEN               => open,                            --                  .arlen
			h2f_ARSIZE              => open,                            --                  .arsize
			h2f_ARBURST             => open,                            --                  .arburst
			h2f_ARLOCK              => open,                            --                  .arlock
			h2f_ARCACHE             => open,                            --                  .arcache
			h2f_ARPROT              => open,                            --                  .arprot
			h2f_ARVALID             => open,                            --                  .arvalid
			h2f_ARREADY             => open,                            --                  .arready
			h2f_RID                 => open,                            --                  .rid
			h2f_RDATA               => open,                            --                  .rdata
			h2f_RRESP               => open,                            --                  .rresp
			h2f_RLAST               => open,                            --                  .rlast
			h2f_RVALID              => open,                            --                  .rvalid
			h2f_RREADY              => open,                            --                  .rready
			f2h_axi_clk             => clk_clk,                         --     f2h_axi_clock.clk
			f2h_AWID                => open,                            --     f2h_axi_slave.awid
			f2h_AWADDR              => open,                            --                  .awaddr
			f2h_AWLEN               => open,                            --                  .awlen
			f2h_AWSIZE              => open,                            --                  .awsize
			f2h_AWBURST             => open,                            --                  .awburst
			f2h_AWLOCK              => open,                            --                  .awlock
			f2h_AWCACHE             => open,                            --                  .awcache
			f2h_AWPROT              => open,                            --                  .awprot
			f2h_AWVALID             => open,                            --                  .awvalid
			f2h_AWREADY             => open,                            --                  .awready
			f2h_AWUSER              => open,                            --                  .awuser
			f2h_WID                 => open,                            --                  .wid
			f2h_WDATA               => open,                            --                  .wdata
			f2h_WSTRB               => open,                            --                  .wstrb
			f2h_WLAST               => open,                            --                  .wlast
			f2h_WVALID              => open,                            --                  .wvalid
			f2h_WREADY              => open,                            --                  .wready
			f2h_BID                 => open,                            --                  .bid
			f2h_BRESP               => open,                            --                  .bresp
			f2h_BVALID              => open,                            --                  .bvalid
			f2h_BREADY              => open,                            --                  .bready
			f2h_ARID                => open,                            --                  .arid
			f2h_ARADDR              => open,                            --                  .araddr
			f2h_ARLEN               => open,                            --                  .arlen
			f2h_ARSIZE              => open,                            --                  .arsize
			f2h_ARBURST             => open,                            --                  .arburst
			f2h_ARLOCK              => open,                            --                  .arlock
			f2h_ARCACHE             => open,                            --                  .arcache
			f2h_ARPROT              => open,                            --                  .arprot
			f2h_ARVALID             => open,                            --                  .arvalid
			f2h_ARREADY             => open,                            --                  .arready
			f2h_ARUSER              => open,                            --                  .aruser
			f2h_RID                 => open,                            --                  .rid
			f2h_RDATA               => open,                            --                  .rdata
			f2h_RRESP               => open,                            --                  .rresp
			f2h_RLAST               => open,                            --                  .rlast
			f2h_RVALID              => open,                            --                  .rvalid
			f2h_RREADY              => open,                            --                  .rready
			h2f_lw_axi_clk          => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID             => open,                            -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR           => open,                            --                  .awaddr
			h2f_lw_AWLEN            => open,                            --                  .awlen
			h2f_lw_AWSIZE           => open,                            --                  .awsize
			h2f_lw_AWBURST          => open,                            --                  .awburst
			h2f_lw_AWLOCK           => open,                            --                  .awlock
			h2f_lw_AWCACHE          => open,                            --                  .awcache
			h2f_lw_AWPROT           => open,                            --                  .awprot
			h2f_lw_AWVALID          => open,                            --                  .awvalid
			h2f_lw_AWREADY          => open,                            --                  .awready
			h2f_lw_WID              => open,                            --                  .wid
			h2f_lw_WDATA            => open,                            --                  .wdata
			h2f_lw_WSTRB            => open,                            --                  .wstrb
			h2f_lw_WLAST            => open,                            --                  .wlast
			h2f_lw_WVALID           => open,                            --                  .wvalid
			h2f_lw_WREADY           => open,                            --                  .wready
			h2f_lw_BID              => open,                            --                  .bid
			h2f_lw_BRESP            => open,                            --                  .bresp
			h2f_lw_BVALID           => open,                            --                  .bvalid
			h2f_lw_BREADY           => open,                            --                  .bready
			h2f_lw_ARID             => open,                            --                  .arid
			h2f_lw_ARADDR           => open,                            --                  .araddr
			h2f_lw_ARLEN            => open,                            --                  .arlen
			h2f_lw_ARSIZE           => open,                            --                  .arsize
			h2f_lw_ARBURST          => open,                            --                  .arburst
			h2f_lw_ARLOCK           => open,                            --                  .arlock
			h2f_lw_ARCACHE          => open,                            --                  .arcache
			h2f_lw_ARPROT           => open,                            --                  .arprot
			h2f_lw_ARVALID          => open,                            --                  .arvalid
			h2f_lw_ARREADY          => open,                            --                  .arready
			h2f_lw_RID              => open,                            --                  .rid
			h2f_lw_RDATA            => open,                            --                  .rdata
			h2f_lw_RRESP            => open,                            --                  .rresp
			h2f_lw_RLAST            => open,                            --                  .rlast
			h2f_lw_RVALID           => open,                            --                  .rvalid
			h2f_lw_RREADY           => open                             --                  .rready
		);

	serial_flash_loader : component altera_serial_flash_loader
		generic map (
			INTENDED_DEVICE_FAMILY  => "Cyclone V",
			ENHANCED_MODE           => true,
			ENABLE_SHARED_ACCESS    => "OFF",
			ENABLE_QUAD_SPI_SUPPORT => true,
			NCSO_WIDTH              => 1
		)
		port map (
			noe_in => serial_flash_loader_0_noe_in_noe  -- noe_in.noe
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	clksampling_clk <= clk_clk;

end architecture rtl; -- of reverbFPGA_Qsys
