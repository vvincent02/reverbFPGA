-- reverbFPGA_Qsys.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity reverbFPGA_Qsys is
	port (
		audio_controller_avalon_left_channel_sink_data     : in    std_logic_vector(23 downto 0) := (others => '0'); --    audio_controller_avalon_left_channel_sink.data
		audio_controller_avalon_left_channel_sink_valid    : in    std_logic                     := '0';             --                                             .valid
		audio_controller_avalon_left_channel_sink_ready    : out   std_logic;                                        --                                             .ready
		audio_controller_avalon_left_channel_source_ready  : in    std_logic                     := '0';             --  audio_controller_avalon_left_channel_source.ready
		audio_controller_avalon_left_channel_source_data   : out   std_logic_vector(23 downto 0);                    --                                             .data
		audio_controller_avalon_left_channel_source_valid  : out   std_logic;                                        --                                             .valid
		audio_controller_avalon_right_channel_sink_data    : in    std_logic_vector(23 downto 0) := (others => '0'); --   audio_controller_avalon_right_channel_sink.data
		audio_controller_avalon_right_channel_sink_valid   : in    std_logic                     := '0';             --                                             .valid
		audio_controller_avalon_right_channel_sink_ready   : out   std_logic;                                        --                                             .ready
		audio_controller_avalon_right_channel_source_ready : in    std_logic                     := '0';             -- audio_controller_avalon_right_channel_source.ready
		audio_controller_avalon_right_channel_source_data  : out   std_logic_vector(23 downto 0);                    --                                             .data
		audio_controller_avalon_right_channel_source_valid : out   std_logic;                                        --                                             .valid
		audio_controller_external_interface_ADCDAT         : in    std_logic                     := '0';             --          audio_controller_external_interface.ADCDAT
		audio_controller_external_interface_ADCLRCK        : in    std_logic                     := '0';             --                                             .ADCLRCK
		audio_controller_external_interface_BCLK           : in    std_logic                     := '0';             --                                             .BCLK
		audio_controller_external_interface_DACDAT         : out   std_logic;                                        --                                             .DACDAT
		audio_controller_external_interface_DACLRCK        : in    std_logic                     := '0';             --                                             .DACLRCK
		audio_pll_0_audio_clk_clk                          : out   std_logic;                                        --                        audio_pll_0_audio_clk.clk
		clk_clk                                            : in    std_logic                     := '0';             --                                          clk.clk
		dampingvalue_pio_external_connection_export        : out   std_logic_vector(24 downto 0);                    --         dampingvalue_pio_external_connection.export
		decayvalue_pio_external_connection_export          : out   std_logic_vector(24 downto 0);                    --           decayvalue_pio_external_connection.export
		hex0_external_connection_export                    : out   std_logic_vector(5 downto 0);                     --                     hex0_external_connection.export
		hex1_external_connection_export                    : out   std_logic_vector(5 downto 0);                     --                     hex1_external_connection.export
		hex2_external_connection_export                    : out   std_logic_vector(5 downto 0);                     --                     hex2_external_connection.export
		hex3_external_connection_export                    : out   std_logic_vector(5 downto 0);                     --                     hex3_external_connection.export
		hex4_external_connection_export                    : out   std_logic_vector(5 downto 0);                     --                     hex4_external_connection.export
		hex5_external_connection_export                    : out   std_logic_vector(5 downto 0);                     --                     hex5_external_connection.export
		hps_io_hps_io_i2c1_inst_SDA                        : inout std_logic                     := '0';             --                                       hps_io.hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL                        : inout std_logic                     := '0';             --                                             .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO48                     : inout std_logic                     := '0';             --                                             .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO53                     : inout std_logic                     := '0';             --                                             .hps_io_gpio_inst_GPIO53
		memory_mem_a                                       : out   std_logic_vector(14 downto 0);                    --                                       memory.mem_a
		memory_mem_ba                                      : out   std_logic_vector(2 downto 0);                     --                                             .mem_ba
		memory_mem_ck                                      : out   std_logic;                                        --                                             .mem_ck
		memory_mem_ck_n                                    : out   std_logic;                                        --                                             .mem_ck_n
		memory_mem_cke                                     : out   std_logic;                                        --                                             .mem_cke
		memory_mem_cs_n                                    : out   std_logic;                                        --                                             .mem_cs_n
		memory_mem_ras_n                                   : out   std_logic;                                        --                                             .mem_ras_n
		memory_mem_cas_n                                   : out   std_logic;                                        --                                             .mem_cas_n
		memory_mem_we_n                                    : out   std_logic;                                        --                                             .mem_we_n
		memory_mem_reset_n                                 : out   std_logic;                                        --                                             .mem_reset_n
		memory_mem_dq                                      : inout std_logic_vector(31 downto 0) := (others => '0'); --                                             .mem_dq
		memory_mem_dqs                                     : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                             .mem_dqs
		memory_mem_dqs_n                                   : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                             .mem_dqs_n
		memory_mem_odt                                     : out   std_logic;                                        --                                             .mem_odt
		memory_mem_dm                                      : out   std_logic_vector(3 downto 0);                     --                                             .mem_dm
		memory_oct_rzqin                                   : in    std_logic                     := '0';             --                                             .oct_rzqin
		mixvalue_pio_external_connection_export            : out   std_logic_vector(23 downto 0);                    --             mixvalue_pio_external_connection.export
		paramtype_pio_external_connection_export           : in    std_logic_vector(3 downto 0)  := (others => '0'); --            paramtype_pio_external_connection.export
		paramvalueupdate_pio_external_connection_export    : in    std_logic_vector(1 downto 0)  := (others => '0'); --     paramvalueupdate_pio_external_connection.export
		predelayvalue_pio_external_connection_export       : out   std_logic_vector(9 downto 0);                     --        predelayvalue_pio_external_connection.export
		reset_reset_n                                      : in    std_logic                     := '0';             --                                        reset.reset_n
		serial_flash_loader_0_noe_in_noe                   : in    std_logic                     := '0'              --                 serial_flash_loader_0_noe_in.noe
	);
end entity reverbFPGA_Qsys;

architecture rtl of reverbFPGA_Qsys is
	component reverbFPGA_Qsys_audio_controller is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset                        : in  std_logic                     := 'X';             -- reset
			from_adc_left_channel_ready  : in  std_logic                     := 'X';             -- ready
			from_adc_left_channel_data   : out std_logic_vector(23 downto 0);                    -- data
			from_adc_left_channel_valid  : out std_logic;                                        -- valid
			from_adc_right_channel_ready : in  std_logic                     := 'X';             -- ready
			from_adc_right_channel_data  : out std_logic_vector(23 downto 0);                    -- data
			from_adc_right_channel_valid : out std_logic;                                        -- valid
			to_dac_left_channel_data     : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_left_channel_valid    : in  std_logic                     := 'X';             -- valid
			to_dac_left_channel_ready    : out std_logic;                                        -- ready
			to_dac_right_channel_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_right_channel_valid   : in  std_logic                     := 'X';             -- valid
			to_dac_right_channel_ready   : out std_logic;                                        -- ready
			AUD_ADCDAT                   : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK                  : in  std_logic                     := 'X';             -- export
			AUD_BCLK                     : in  std_logic                     := 'X';             -- export
			AUD_DACDAT                   : out std_logic;                                        -- export
			AUD_DACLRCK                  : in  std_logic                     := 'X'              -- export
		);
	end component reverbFPGA_Qsys_audio_controller;

	component reverbFPGA_Qsys_audio_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component reverbFPGA_Qsys_audio_pll_0;

	component reverbFPGA_Qsys_dampingValue_PIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(24 downto 0)                     -- export
		);
	end component reverbFPGA_Qsys_dampingValue_PIO;

	component reverbFPGA_Qsys_hex0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(5 downto 0)                      -- export
		);
	end component reverbFPGA_Qsys_hex0;

	component reverbFPGA_Qsys_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                   : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                  : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                  : out   std_logic;                                        -- mem_ck
			mem_ck_n                : out   std_logic;                                        -- mem_ck_n
			mem_cke                 : out   std_logic;                                        -- mem_cke
			mem_cs_n                : out   std_logic;                                        -- mem_cs_n
			mem_ras_n               : out   std_logic;                                        -- mem_ras_n
			mem_cas_n               : out   std_logic;                                        -- mem_cas_n
			mem_we_n                : out   std_logic;                                        -- mem_we_n
			mem_reset_n             : out   std_logic;                                        -- mem_reset_n
			mem_dq                  : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                 : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n               : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                 : out   std_logic;                                        -- mem_odt
			mem_dm                  : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin               : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_i2c1_inst_SDA    : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL    : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO48 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			h2f_rst_n               : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk          : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID             : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR           : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN            : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE           : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST          : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK           : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE          : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT           : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID          : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY          : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID              : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA            : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB            : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST            : out   std_logic;                                        -- wlast
			h2f_lw_WVALID           : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY           : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID              : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP            : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID           : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY           : out   std_logic;                                        -- bready
			h2f_lw_ARID             : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR           : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN            : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE           : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST          : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK           : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE          : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT           : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID          : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY          : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID              : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA            : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP            : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST            : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID           : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY           : out   std_logic                                         -- rready
		);
	end component reverbFPGA_Qsys_hps_0;

	component reverbFPGA_Qsys_mixValue_PIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(23 downto 0)                     -- export
		);
	end component reverbFPGA_Qsys_mixValue_PIO;

	component reverbFPGA_Qsys_paramType_PIO is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component reverbFPGA_Qsys_paramType_PIO;

	component reverbFPGA_Qsys_paramValueUpdate_PIO is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component reverbFPGA_Qsys_paramValueUpdate_PIO;

	component reverbFPGA_Qsys_preDelayValue_PIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component reverbFPGA_Qsys_preDelayValue_PIO;

	component altera_serial_flash_loader is
		generic (
			INTENDED_DEVICE_FAMILY  : string  := "";
			ENHANCED_MODE           : boolean := true;
			ENABLE_SHARED_ACCESS    : string  := "OFF";
			ENABLE_QUAD_SPI_SUPPORT : boolean := false;
			NCSO_WIDTH              : integer := 1
		);
		port (
			noe_in : in std_logic := 'X'  -- noe
		);
	end component altera_serial_flash_loader;

	component reverbFPGA_Qsys_mm_interconnect_0 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			dampingValue_PIO_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			dampingValue_PIO_s1_address                                         : out std_logic_vector(1 downto 0);                     -- address
			dampingValue_PIO_s1_write                                           : out std_logic;                                        -- write
			dampingValue_PIO_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dampingValue_PIO_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			dampingValue_PIO_s1_chipselect                                      : out std_logic;                                        -- chipselect
			decayValue_PIO_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			decayValue_PIO_s1_write                                             : out std_logic;                                        -- write
			decayValue_PIO_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			decayValue_PIO_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			decayValue_PIO_s1_chipselect                                        : out std_logic;                                        -- chipselect
			hex0_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			hex0_s1_write                                                       : out std_logic;                                        -- write
			hex0_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex0_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			hex0_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			hex1_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			hex1_s1_write                                                       : out std_logic;                                        -- write
			hex1_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex1_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			hex1_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			hex2_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			hex2_s1_write                                                       : out std_logic;                                        -- write
			hex2_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex2_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			hex2_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			hex3_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			hex3_s1_write                                                       : out std_logic;                                        -- write
			hex3_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex3_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			hex3_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			hex4_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			hex4_s1_write                                                       : out std_logic;                                        -- write
			hex4_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex4_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			hex4_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			hex5_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			hex5_s1_write                                                       : out std_logic;                                        -- write
			hex5_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex5_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			hex5_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			mixValue_PIO_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			mixValue_PIO_s1_write                                               : out std_logic;                                        -- write
			mixValue_PIO_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mixValue_PIO_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			mixValue_PIO_s1_chipselect                                          : out std_logic;                                        -- chipselect
			paramType_PIO_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			paramType_PIO_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			paramValueUpdate_PIO_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			paramValueUpdate_PIO_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			preDelayValue_PIO_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			preDelayValue_PIO_s1_write                                          : out std_logic;                                        -- write
			preDelayValue_PIO_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			preDelayValue_PIO_s1_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			preDelayValue_PIO_s1_chipselect                                     : out std_logic                                         -- chipselect
		);
	end component reverbFPGA_Qsys_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal hps_0_h2f_lw_axi_master_awburst                        : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                          : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                          : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                         : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                            : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                         : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                          : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                            : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                        : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                         : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                         : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                         : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                         : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                          : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                        : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                        : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                           : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                         : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                         : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                         : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                        : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                        : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                        : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                         : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                         : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                          : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                          : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                           : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                            : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                         : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                         : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                        : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                         : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_0_dampingvalue_pio_s1_chipselect       : std_logic;                     -- mm_interconnect_0:dampingValue_PIO_s1_chipselect -> dampingValue_PIO:chipselect
	signal mm_interconnect_0_dampingvalue_pio_s1_readdata         : std_logic_vector(31 downto 0); -- dampingValue_PIO:readdata -> mm_interconnect_0:dampingValue_PIO_s1_readdata
	signal mm_interconnect_0_dampingvalue_pio_s1_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:dampingValue_PIO_s1_address -> dampingValue_PIO:address
	signal mm_interconnect_0_dampingvalue_pio_s1_write            : std_logic;                     -- mm_interconnect_0:dampingValue_PIO_s1_write -> mm_interconnect_0_dampingvalue_pio_s1_write:in
	signal mm_interconnect_0_dampingvalue_pio_s1_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:dampingValue_PIO_s1_writedata -> dampingValue_PIO:writedata
	signal mm_interconnect_0_mixvalue_pio_s1_chipselect           : std_logic;                     -- mm_interconnect_0:mixValue_PIO_s1_chipselect -> mixValue_PIO:chipselect
	signal mm_interconnect_0_mixvalue_pio_s1_readdata             : std_logic_vector(31 downto 0); -- mixValue_PIO:readdata -> mm_interconnect_0:mixValue_PIO_s1_readdata
	signal mm_interconnect_0_mixvalue_pio_s1_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mixValue_PIO_s1_address -> mixValue_PIO:address
	signal mm_interconnect_0_mixvalue_pio_s1_write                : std_logic;                     -- mm_interconnect_0:mixValue_PIO_s1_write -> mm_interconnect_0_mixvalue_pio_s1_write:in
	signal mm_interconnect_0_mixvalue_pio_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:mixValue_PIO_s1_writedata -> mixValue_PIO:writedata
	signal mm_interconnect_0_paramvalueupdate_pio_s1_readdata     : std_logic_vector(31 downto 0); -- paramValueUpdate_PIO:readdata -> mm_interconnect_0:paramValueUpdate_PIO_s1_readdata
	signal mm_interconnect_0_paramvalueupdate_pio_s1_address      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:paramValueUpdate_PIO_s1_address -> paramValueUpdate_PIO:address
	signal mm_interconnect_0_paramtype_pio_s1_readdata            : std_logic_vector(31 downto 0); -- paramType_PIO:readdata -> mm_interconnect_0:paramType_PIO_s1_readdata
	signal mm_interconnect_0_paramtype_pio_s1_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:paramType_PIO_s1_address -> paramType_PIO:address
	signal mm_interconnect_0_decayvalue_pio_s1_chipselect         : std_logic;                     -- mm_interconnect_0:decayValue_PIO_s1_chipselect -> decayValue_PIO:chipselect
	signal mm_interconnect_0_decayvalue_pio_s1_readdata           : std_logic_vector(31 downto 0); -- decayValue_PIO:readdata -> mm_interconnect_0:decayValue_PIO_s1_readdata
	signal mm_interconnect_0_decayvalue_pio_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:decayValue_PIO_s1_address -> decayValue_PIO:address
	signal mm_interconnect_0_decayvalue_pio_s1_write              : std_logic;                     -- mm_interconnect_0:decayValue_PIO_s1_write -> mm_interconnect_0_decayvalue_pio_s1_write:in
	signal mm_interconnect_0_decayvalue_pio_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:decayValue_PIO_s1_writedata -> decayValue_PIO:writedata
	signal mm_interconnect_0_hex0_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:hex0_s1_chipselect -> hex0:chipselect
	signal mm_interconnect_0_hex0_s1_readdata                     : std_logic_vector(31 downto 0); -- hex0:readdata -> mm_interconnect_0:hex0_s1_readdata
	signal mm_interconnect_0_hex0_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex0_s1_address -> hex0:address
	signal mm_interconnect_0_hex0_s1_write                        : std_logic;                     -- mm_interconnect_0:hex0_s1_write -> mm_interconnect_0_hex0_s1_write:in
	signal mm_interconnect_0_hex0_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex0_s1_writedata -> hex0:writedata
	signal mm_interconnect_0_hex1_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:hex1_s1_chipselect -> hex1:chipselect
	signal mm_interconnect_0_hex1_s1_readdata                     : std_logic_vector(31 downto 0); -- hex1:readdata -> mm_interconnect_0:hex1_s1_readdata
	signal mm_interconnect_0_hex1_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex1_s1_address -> hex1:address
	signal mm_interconnect_0_hex1_s1_write                        : std_logic;                     -- mm_interconnect_0:hex1_s1_write -> mm_interconnect_0_hex1_s1_write:in
	signal mm_interconnect_0_hex1_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex1_s1_writedata -> hex1:writedata
	signal mm_interconnect_0_hex2_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:hex2_s1_chipselect -> hex2:chipselect
	signal mm_interconnect_0_hex2_s1_readdata                     : std_logic_vector(31 downto 0); -- hex2:readdata -> mm_interconnect_0:hex2_s1_readdata
	signal mm_interconnect_0_hex2_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex2_s1_address -> hex2:address
	signal mm_interconnect_0_hex2_s1_write                        : std_logic;                     -- mm_interconnect_0:hex2_s1_write -> mm_interconnect_0_hex2_s1_write:in
	signal mm_interconnect_0_hex2_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex2_s1_writedata -> hex2:writedata
	signal mm_interconnect_0_hex3_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:hex3_s1_chipselect -> hex3:chipselect
	signal mm_interconnect_0_hex3_s1_readdata                     : std_logic_vector(31 downto 0); -- hex3:readdata -> mm_interconnect_0:hex3_s1_readdata
	signal mm_interconnect_0_hex3_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex3_s1_address -> hex3:address
	signal mm_interconnect_0_hex3_s1_write                        : std_logic;                     -- mm_interconnect_0:hex3_s1_write -> mm_interconnect_0_hex3_s1_write:in
	signal mm_interconnect_0_hex3_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex3_s1_writedata -> hex3:writedata
	signal mm_interconnect_0_hex4_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:hex4_s1_chipselect -> hex4:chipselect
	signal mm_interconnect_0_hex4_s1_readdata                     : std_logic_vector(31 downto 0); -- hex4:readdata -> mm_interconnect_0:hex4_s1_readdata
	signal mm_interconnect_0_hex4_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex4_s1_address -> hex4:address
	signal mm_interconnect_0_hex4_s1_write                        : std_logic;                     -- mm_interconnect_0:hex4_s1_write -> mm_interconnect_0_hex4_s1_write:in
	signal mm_interconnect_0_hex4_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex4_s1_writedata -> hex4:writedata
	signal mm_interconnect_0_hex5_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:hex5_s1_chipselect -> hex5:chipselect
	signal mm_interconnect_0_hex5_s1_readdata                     : std_logic_vector(31 downto 0); -- hex5:readdata -> mm_interconnect_0:hex5_s1_readdata
	signal mm_interconnect_0_hex5_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex5_s1_address -> hex5:address
	signal mm_interconnect_0_hex5_s1_write                        : std_logic;                     -- mm_interconnect_0:hex5_s1_write -> mm_interconnect_0_hex5_s1_write:in
	signal mm_interconnect_0_hex5_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex5_s1_writedata -> hex5:writedata
	signal mm_interconnect_0_predelayvalue_pio_s1_chipselect      : std_logic;                     -- mm_interconnect_0:preDelayValue_PIO_s1_chipselect -> preDelayValue_PIO:chipselect
	signal mm_interconnect_0_predelayvalue_pio_s1_readdata        : std_logic_vector(31 downto 0); -- preDelayValue_PIO:readdata -> mm_interconnect_0:preDelayValue_PIO_s1_readdata
	signal mm_interconnect_0_predelayvalue_pio_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:preDelayValue_PIO_s1_address -> preDelayValue_PIO:address
	signal mm_interconnect_0_predelayvalue_pio_s1_write           : std_logic;                     -- mm_interconnect_0:preDelayValue_PIO_s1_write -> mm_interconnect_0_predelayvalue_pio_s1_write:in
	signal mm_interconnect_0_predelayvalue_pio_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:preDelayValue_PIO_s1_writedata -> preDelayValue_PIO:writedata
	signal rst_controller_reset_out_reset                         : std_logic;                     -- rst_controller:reset_out -> [audio_controller:reset, mm_interconnect_0:dampingValue_PIO_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                     : std_logic;                     -- rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal hps_0_h2f_reset_reset                                  : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal reset_reset_n_ports_inv                                : std_logic;                     -- reset_reset_n:inv -> [audio_pll_0:ref_reset_reset, rst_controller:reset_in0]
	signal mm_interconnect_0_dampingvalue_pio_s1_write_ports_inv  : std_logic;                     -- mm_interconnect_0_dampingvalue_pio_s1_write:inv -> dampingValue_PIO:write_n
	signal mm_interconnect_0_mixvalue_pio_s1_write_ports_inv      : std_logic;                     -- mm_interconnect_0_mixvalue_pio_s1_write:inv -> mixValue_PIO:write_n
	signal mm_interconnect_0_decayvalue_pio_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_decayvalue_pio_s1_write:inv -> decayValue_PIO:write_n
	signal mm_interconnect_0_hex0_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_hex0_s1_write:inv -> hex0:write_n
	signal mm_interconnect_0_hex1_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_hex1_s1_write:inv -> hex1:write_n
	signal mm_interconnect_0_hex2_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_hex2_s1_write:inv -> hex2:write_n
	signal mm_interconnect_0_hex3_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_hex3_s1_write:inv -> hex3:write_n
	signal mm_interconnect_0_hex4_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_hex4_s1_write:inv -> hex4:write_n
	signal mm_interconnect_0_hex5_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_hex5_s1_write:inv -> hex5:write_n
	signal mm_interconnect_0_predelayvalue_pio_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_predelayvalue_pio_s1_write:inv -> preDelayValue_PIO:write_n
	signal rst_controller_reset_out_reset_ports_inv               : std_logic;                     -- rst_controller_reset_out_reset:inv -> [dampingValue_PIO:reset_n, decayValue_PIO:reset_n, hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, mixValue_PIO:reset_n, paramType_PIO:reset_n, paramValueUpdate_PIO:reset_n, preDelayValue_PIO:reset_n]
	signal hps_0_h2f_reset_reset_ports_inv                        : std_logic;                     -- hps_0_h2f_reset_reset:inv -> rst_controller_001:reset_in0

begin

	audio_controller : component reverbFPGA_Qsys_audio_controller
		port map (
			clk                          => clk_clk,                                            --                         clk.clk
			reset                        => rst_controller_reset_out_reset,                     --                       reset.reset
			from_adc_left_channel_ready  => audio_controller_avalon_left_channel_source_ready,  --  avalon_left_channel_source.ready
			from_adc_left_channel_data   => audio_controller_avalon_left_channel_source_data,   --                            .data
			from_adc_left_channel_valid  => audio_controller_avalon_left_channel_source_valid,  --                            .valid
			from_adc_right_channel_ready => audio_controller_avalon_right_channel_source_ready, -- avalon_right_channel_source.ready
			from_adc_right_channel_data  => audio_controller_avalon_right_channel_source_data,  --                            .data
			from_adc_right_channel_valid => audio_controller_avalon_right_channel_source_valid, --                            .valid
			to_dac_left_channel_data     => audio_controller_avalon_left_channel_sink_data,     --    avalon_left_channel_sink.data
			to_dac_left_channel_valid    => audio_controller_avalon_left_channel_sink_valid,    --                            .valid
			to_dac_left_channel_ready    => audio_controller_avalon_left_channel_sink_ready,    --                            .ready
			to_dac_right_channel_data    => audio_controller_avalon_right_channel_sink_data,    --   avalon_right_channel_sink.data
			to_dac_right_channel_valid   => audio_controller_avalon_right_channel_sink_valid,   --                            .valid
			to_dac_right_channel_ready   => audio_controller_avalon_right_channel_sink_ready,   --                            .ready
			AUD_ADCDAT                   => audio_controller_external_interface_ADCDAT,         --          external_interface.export
			AUD_ADCLRCK                  => audio_controller_external_interface_ADCLRCK,        --                            .export
			AUD_BCLK                     => audio_controller_external_interface_BCLK,           --                            .export
			AUD_DACDAT                   => audio_controller_external_interface_DACDAT,         --                            .export
			AUD_DACLRCK                  => audio_controller_external_interface_DACLRCK         --                            .export
		);

	audio_pll_0 : component reverbFPGA_Qsys_audio_pll_0
		port map (
			ref_clk_clk        => clk_clk,                   --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,   --    ref_reset.reset
			audio_clk_clk      => audio_pll_0_audio_clk_clk, --    audio_clk.clk
			reset_source_reset => open                       -- reset_source.reset
		);

	dampingvalue_pio : component reverbFPGA_Qsys_dampingValue_PIO
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_dampingvalue_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_dampingvalue_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_dampingvalue_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_dampingvalue_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_dampingvalue_pio_s1_readdata,        --                    .readdata
			out_port   => dampingvalue_pio_external_connection_export            -- external_connection.export
		);

	decayvalue_pio : component reverbFPGA_Qsys_dampingValue_PIO
		port map (
			clk        => clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => mm_interconnect_0_decayvalue_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_decayvalue_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_decayvalue_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_decayvalue_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_decayvalue_pio_s1_readdata,        --                    .readdata
			out_port   => decayvalue_pio_external_connection_export            -- external_connection.export
		);

	hex0 : component reverbFPGA_Qsys_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex0_s1_readdata,        --                    .readdata
			out_port   => hex0_external_connection_export            -- external_connection.export
		);

	hex1 : component reverbFPGA_Qsys_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex1_s1_readdata,        --                    .readdata
			out_port   => hex1_external_connection_export            -- external_connection.export
		);

	hex2 : component reverbFPGA_Qsys_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex2_s1_readdata,        --                    .readdata
			out_port   => hex2_external_connection_export            -- external_connection.export
		);

	hex3 : component reverbFPGA_Qsys_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex3_s1_readdata,        --                    .readdata
			out_port   => hex3_external_connection_export            -- external_connection.export
		);

	hex4 : component reverbFPGA_Qsys_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex4_s1_readdata,        --                    .readdata
			out_port   => hex4_external_connection_export            -- external_connection.export
		);

	hex5 : component reverbFPGA_Qsys_hex0
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_hex5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex5_s1_readdata,        --                    .readdata
			out_port   => hex5_external_connection_export            -- external_connection.export
		);

	hps_0 : component reverbFPGA_Qsys_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                   => memory_mem_a,                    --            memory.mem_a
			mem_ba                  => memory_mem_ba,                   --                  .mem_ba
			mem_ck                  => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n                => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                 => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n                => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n               => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n               => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n             => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq                  => memory_mem_dq,                   --                  .mem_dq
			mem_dqs                 => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n               => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                 => memory_mem_odt,                  --                  .mem_odt
			mem_dm                  => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin               => memory_oct_rzqin,                --                  .oct_rzqin
			hps_io_i2c1_inst_SDA    => hps_io_hps_io_i2c1_inst_SDA,     --            hps_io.hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL    => hps_io_hps_io_i2c1_inst_SCL,     --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO48 => hps_io_hps_io_gpio_inst_GPIO48,  --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53 => hps_io_hps_io_gpio_inst_GPIO53,  --                  .hps_io_gpio_inst_GPIO53
			h2f_rst_n               => hps_0_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_lw_axi_clk          => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID             => hps_0_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR           => hps_0_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN            => hps_0_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE           => hps_0_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST          => hps_0_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK           => hps_0_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE          => hps_0_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT           => hps_0_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID          => hps_0_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY          => hps_0_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID              => hps_0_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA            => hps_0_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB            => hps_0_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST            => hps_0_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID           => hps_0_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY           => hps_0_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID              => hps_0_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP            => hps_0_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID           => hps_0_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY           => hps_0_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID             => hps_0_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR           => hps_0_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN            => hps_0_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE           => hps_0_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST          => hps_0_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK           => hps_0_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE          => hps_0_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT           => hps_0_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID          => hps_0_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY          => hps_0_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID              => hps_0_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA            => hps_0_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP            => hps_0_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST            => hps_0_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID           => hps_0_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY           => hps_0_h2f_lw_axi_master_rready   --                  .rready
		);

	mixvalue_pio : component reverbFPGA_Qsys_mixValue_PIO
		port map (
			clk        => clk_clk,                                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_mixvalue_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_mixvalue_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_mixvalue_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_mixvalue_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_mixvalue_pio_s1_readdata,        --                    .readdata
			out_port   => mixvalue_pio_external_connection_export            -- external_connection.export
		);

	paramtype_pio : component reverbFPGA_Qsys_paramType_PIO
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => mm_interconnect_0_paramtype_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_paramtype_pio_s1_readdata, --                    .readdata
			in_port  => paramtype_pio_external_connection_export     -- external_connection.export
		);

	paramvalueupdate_pio : component reverbFPGA_Qsys_paramValueUpdate_PIO
		port map (
			clk      => clk_clk,                                            --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address  => mm_interconnect_0_paramvalueupdate_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_paramvalueupdate_pio_s1_readdata, --                    .readdata
			in_port  => paramvalueupdate_pio_external_connection_export     -- external_connection.export
		);

	predelayvalue_pio : component reverbFPGA_Qsys_preDelayValue_PIO
		port map (
			clk        => clk_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,               --               reset.reset_n
			address    => mm_interconnect_0_predelayvalue_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_predelayvalue_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_predelayvalue_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_predelayvalue_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_predelayvalue_pio_s1_readdata,        --                    .readdata
			out_port   => predelayvalue_pio_external_connection_export            -- external_connection.export
		);

	serial_flash_loader : component altera_serial_flash_loader
		generic map (
			INTENDED_DEVICE_FAMILY  => "Cyclone V",
			ENHANCED_MODE           => true,
			ENABLE_SHARED_ACCESS    => "OFF",
			ENABLE_QUAD_SPI_SUPPORT => true,
			NCSO_WIDTH              => 1
		)
		port map (
			noe_in => serial_flash_loader_0_noe_in_noe  -- noe_in.noe
		);

	mm_interconnect_0 : component reverbFPGA_Qsys_mm_interconnect_0
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                       --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                     --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                      --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                     --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                    --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                     --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                    --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                     --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                    --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                    --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                        --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                      --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                      --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                      --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                     --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                     --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                        --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                      --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                     --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                     --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                       --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                     --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                      --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                     --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                    --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                     --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                    --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                     --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                    --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                    --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                        --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                      --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                      --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                      --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                     --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                     --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                            --                                                     clk_0_clk.clk
			dampingValue_PIO_reset_reset_bridge_in_reset_reset                  => rst_controller_reset_out_reset,                     --                  dampingValue_PIO_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                 -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			dampingValue_PIO_s1_address                                         => mm_interconnect_0_dampingvalue_pio_s1_address,      --                                           dampingValue_PIO_s1.address
			dampingValue_PIO_s1_write                                           => mm_interconnect_0_dampingvalue_pio_s1_write,        --                                                              .write
			dampingValue_PIO_s1_readdata                                        => mm_interconnect_0_dampingvalue_pio_s1_readdata,     --                                                              .readdata
			dampingValue_PIO_s1_writedata                                       => mm_interconnect_0_dampingvalue_pio_s1_writedata,    --                                                              .writedata
			dampingValue_PIO_s1_chipselect                                      => mm_interconnect_0_dampingvalue_pio_s1_chipselect,   --                                                              .chipselect
			decayValue_PIO_s1_address                                           => mm_interconnect_0_decayvalue_pio_s1_address,        --                                             decayValue_PIO_s1.address
			decayValue_PIO_s1_write                                             => mm_interconnect_0_decayvalue_pio_s1_write,          --                                                              .write
			decayValue_PIO_s1_readdata                                          => mm_interconnect_0_decayvalue_pio_s1_readdata,       --                                                              .readdata
			decayValue_PIO_s1_writedata                                         => mm_interconnect_0_decayvalue_pio_s1_writedata,      --                                                              .writedata
			decayValue_PIO_s1_chipselect                                        => mm_interconnect_0_decayvalue_pio_s1_chipselect,     --                                                              .chipselect
			hex0_s1_address                                                     => mm_interconnect_0_hex0_s1_address,                  --                                                       hex0_s1.address
			hex0_s1_write                                                       => mm_interconnect_0_hex0_s1_write,                    --                                                              .write
			hex0_s1_readdata                                                    => mm_interconnect_0_hex0_s1_readdata,                 --                                                              .readdata
			hex0_s1_writedata                                                   => mm_interconnect_0_hex0_s1_writedata,                --                                                              .writedata
			hex0_s1_chipselect                                                  => mm_interconnect_0_hex0_s1_chipselect,               --                                                              .chipselect
			hex1_s1_address                                                     => mm_interconnect_0_hex1_s1_address,                  --                                                       hex1_s1.address
			hex1_s1_write                                                       => mm_interconnect_0_hex1_s1_write,                    --                                                              .write
			hex1_s1_readdata                                                    => mm_interconnect_0_hex1_s1_readdata,                 --                                                              .readdata
			hex1_s1_writedata                                                   => mm_interconnect_0_hex1_s1_writedata,                --                                                              .writedata
			hex1_s1_chipselect                                                  => mm_interconnect_0_hex1_s1_chipselect,               --                                                              .chipselect
			hex2_s1_address                                                     => mm_interconnect_0_hex2_s1_address,                  --                                                       hex2_s1.address
			hex2_s1_write                                                       => mm_interconnect_0_hex2_s1_write,                    --                                                              .write
			hex2_s1_readdata                                                    => mm_interconnect_0_hex2_s1_readdata,                 --                                                              .readdata
			hex2_s1_writedata                                                   => mm_interconnect_0_hex2_s1_writedata,                --                                                              .writedata
			hex2_s1_chipselect                                                  => mm_interconnect_0_hex2_s1_chipselect,               --                                                              .chipselect
			hex3_s1_address                                                     => mm_interconnect_0_hex3_s1_address,                  --                                                       hex3_s1.address
			hex3_s1_write                                                       => mm_interconnect_0_hex3_s1_write,                    --                                                              .write
			hex3_s1_readdata                                                    => mm_interconnect_0_hex3_s1_readdata,                 --                                                              .readdata
			hex3_s1_writedata                                                   => mm_interconnect_0_hex3_s1_writedata,                --                                                              .writedata
			hex3_s1_chipselect                                                  => mm_interconnect_0_hex3_s1_chipselect,               --                                                              .chipselect
			hex4_s1_address                                                     => mm_interconnect_0_hex4_s1_address,                  --                                                       hex4_s1.address
			hex4_s1_write                                                       => mm_interconnect_0_hex4_s1_write,                    --                                                              .write
			hex4_s1_readdata                                                    => mm_interconnect_0_hex4_s1_readdata,                 --                                                              .readdata
			hex4_s1_writedata                                                   => mm_interconnect_0_hex4_s1_writedata,                --                                                              .writedata
			hex4_s1_chipselect                                                  => mm_interconnect_0_hex4_s1_chipselect,               --                                                              .chipselect
			hex5_s1_address                                                     => mm_interconnect_0_hex5_s1_address,                  --                                                       hex5_s1.address
			hex5_s1_write                                                       => mm_interconnect_0_hex5_s1_write,                    --                                                              .write
			hex5_s1_readdata                                                    => mm_interconnect_0_hex5_s1_readdata,                 --                                                              .readdata
			hex5_s1_writedata                                                   => mm_interconnect_0_hex5_s1_writedata,                --                                                              .writedata
			hex5_s1_chipselect                                                  => mm_interconnect_0_hex5_s1_chipselect,               --                                                              .chipselect
			mixValue_PIO_s1_address                                             => mm_interconnect_0_mixvalue_pio_s1_address,          --                                               mixValue_PIO_s1.address
			mixValue_PIO_s1_write                                               => mm_interconnect_0_mixvalue_pio_s1_write,            --                                                              .write
			mixValue_PIO_s1_readdata                                            => mm_interconnect_0_mixvalue_pio_s1_readdata,         --                                                              .readdata
			mixValue_PIO_s1_writedata                                           => mm_interconnect_0_mixvalue_pio_s1_writedata,        --                                                              .writedata
			mixValue_PIO_s1_chipselect                                          => mm_interconnect_0_mixvalue_pio_s1_chipselect,       --                                                              .chipselect
			paramType_PIO_s1_address                                            => mm_interconnect_0_paramtype_pio_s1_address,         --                                              paramType_PIO_s1.address
			paramType_PIO_s1_readdata                                           => mm_interconnect_0_paramtype_pio_s1_readdata,        --                                                              .readdata
			paramValueUpdate_PIO_s1_address                                     => mm_interconnect_0_paramvalueupdate_pio_s1_address,  --                                       paramValueUpdate_PIO_s1.address
			paramValueUpdate_PIO_s1_readdata                                    => mm_interconnect_0_paramvalueupdate_pio_s1_readdata, --                                                              .readdata
			preDelayValue_PIO_s1_address                                        => mm_interconnect_0_predelayvalue_pio_s1_address,     --                                          preDelayValue_PIO_s1.address
			preDelayValue_PIO_s1_write                                          => mm_interconnect_0_predelayvalue_pio_s1_write,       --                                                              .write
			preDelayValue_PIO_s1_readdata                                       => mm_interconnect_0_predelayvalue_pio_s1_readdata,    --                                                              .readdata
			preDelayValue_PIO_s1_writedata                                      => mm_interconnect_0_predelayvalue_pio_s1_writedata,   --                                                              .writedata
			preDelayValue_PIO_s1_chipselect                                     => mm_interconnect_0_predelayvalue_pio_s1_chipselect   --                                                              .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_dampingvalue_pio_s1_write_ports_inv <= not mm_interconnect_0_dampingvalue_pio_s1_write;

	mm_interconnect_0_mixvalue_pio_s1_write_ports_inv <= not mm_interconnect_0_mixvalue_pio_s1_write;

	mm_interconnect_0_decayvalue_pio_s1_write_ports_inv <= not mm_interconnect_0_decayvalue_pio_s1_write;

	mm_interconnect_0_hex0_s1_write_ports_inv <= not mm_interconnect_0_hex0_s1_write;

	mm_interconnect_0_hex1_s1_write_ports_inv <= not mm_interconnect_0_hex1_s1_write;

	mm_interconnect_0_hex2_s1_write_ports_inv <= not mm_interconnect_0_hex2_s1_write;

	mm_interconnect_0_hex3_s1_write_ports_inv <= not mm_interconnect_0_hex3_s1_write;

	mm_interconnect_0_hex4_s1_write_ports_inv <= not mm_interconnect_0_hex4_s1_write;

	mm_interconnect_0_hex5_s1_write_ports_inv <= not mm_interconnect_0_hex5_s1_write;

	mm_interconnect_0_predelayvalue_pio_s1_write_ports_inv <= not mm_interconnect_0_predelayvalue_pio_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of reverbFPGA_Qsys
